LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.conv_integer;

ENTITY InstructionMemory IS PORT (
    addr : IN std_logic_vector(7 DOWNTO 0);
    data : OUT std_logic_vector(31 DOWNTO 0));
END ENTITY;

ARCHITECTURE Behavioral OF InstructionMemory IS
    TYPE mem_t IS ARRAY (0 TO 255) OF std_logic_vector(31 DOWNTO 0);

    CONSTANT switch_chanel : mem_t := (
    x"14010000", --read r1 1
    x"14020100", --read r2 2 
    x"0C000101", --print r1 2
    x"0C000002", --print r2 1
    x"07000000", --jump 0
    OTHERS => (OTHERS => '0'));

    CONSTANT papa_noel : mem_t := (
    x"06020200", -- 00# afc r2 2
    x"06010100", -- 01# afc r1 1
    x"06000100", -- 02# afc r0 1
    x"08000200", -- 03# jmf 2 r0 
    x"06057F00", -- 04# afc r5 7F
    x"06047F00", -- 05# afc r4 7F
    x"06037F00", -- 06# afc r3 7F
    x"03030301", -- 07# sub r3 r3 r1
    x"08000A03", -- 08# jmf A r3
    x"07000700", -- 09# jmp 7
    x"03040401", -- 0A# sub r4 r4 r1
    x"08000D04", -- 0B# jmf D r4
    x"07000600", -- 0C# jmp 6
    x"03050501", -- 0D# sub r5 r5 r1
    x"08001005", -- 0E# jmf 10 r5
    x"07000500", -- 0F# jmp 5
    x"0C000000", -- 10# print r0 1
    x"0C000100", -- 11# print r0 2
    x"02000002", -- 12# mul r0 r0 r2
    x"07000300", -- 13# jmp 3
    OTHERS => (OTHERS => '0'));

    CONSTANT program1 : mem_t := (-- marche pas :c
    x"06010200",
    x"01000001",
    x"07000400",
    x"00000000",
    x"06010100",
    x"06020000",
    x"01020200",
    x"11000102",
    x"06010000",
    x"01010100",
    x"10010001",
    x"08001D01",
    x"14010100",
    x"06020000",
    x"01020200",
    x"11000102",
    x"06010000",
    x"01010100",
    x"10010001",
    x"0C000001",
    x"14010000",
    x"06020000",
    x"01020200",
    x"11000102",
    x"06010000",
    x"01010100",
    x"10010001",
    x"0C000101",
    x"07000400",
    OTHERS => (OTHERS => '0'));

    CONSTANT program2 : mem_t := (-- marche pas :c
    x"06010100",
    x"01000001",
    x"07000300",
    x"06010000",
    x"06020000",
    x"01020200",
    x"11000102",
    x"06010000",
    x"06020100",
    x"01020200",
    x"11000102",
    x"06010100",
    x"01010100",
    x"10010001",
    x"06020000",
    x"01020200",
    x"11000102",
    x"06010100",
    x"06020100",
    x"01020200",
    x"11000102",
    x"06010100",
    x"01010100",
    x"10010001",
    x"0800C701",
    x"06010000",
    x"06020100",
    x"01020200",
    x"11000102",
    x"06020100",
    x"01020200",
    x"10020002",
    x"06010000",
    x"01010100",
    x"10010001",
    x"0B010102",
    x"06020100",
    x"01020200",
    x"11000102",
    x"06010100",
    x"01010100",
    x"10010001",
    x"08003501",
    x"06010100",
    x"06020100",
    x"01020200",
    x"11000102",
    x"06010100",
    x"01010100",
    x"10010001",
    x"06020000",
    x"01020200",
    x"11000102",
    x"06010000",
    x"06020100",
    x"01020200",
    x"11000102",
    x"06011000",
    x"06020200",
    x"01020200",
    x"11000102",
    x"06010200",
    x"01010100",
    x"10010001",
    x"06020100",
    x"01020200",
    x"11000102",
    x"06010100",
    x"01010100",
    x"10010001",
    x"0800AA01",
    x"06010100",
    x"06020200",
    x"01020200",
    x"11000102",
    x"06020200",
    x"01020200",
    x"10020002",
    x"06010100",
    x"01010100",
    x"10010001",
    x"03010102",
    x"06020200",
    x"01020200",
    x"11000102",
    x"06010200",
    x"01010100",
    x"10010001",
    x"06020100",
    x"01020200",
    x"11000102",
    x"06010000",
    x"06020200",
    x"01020200",
    x"11000102",
    x"06011000",
    x"06020300",
    x"01020200",
    x"11000102",
    x"06010300",
    x"01010100",
    x"10010001",
    x"06020200",
    x"01020200",
    x"11000102",
    x"06010200",
    x"01010100",
    x"10010001",
    x"0800A901",
    x"06010100",
    x"06020300",
    x"01020200",
    x"11000102",
    x"06020300",
    x"01020200",
    x"10020002",
    x"06010200",
    x"01010100",
    x"10010001",
    x"03010102",
    x"06020300",
    x"01020200",
    x"11000102",
    x"06010300",
    x"01010100",
    x"10010001",
    x"06020200",
    x"01020200",
    x"11000102",
    x"06010000",
    x"06020300",
    x"01020200",
    x"11000102",
    x"06011000",
    x"06020400",
    x"01020200",
    x"11000102",
    x"06010400",
    x"01010100",
    x"10010001",
    x"06020300",
    x"01020200",
    x"11000102",
    x"06010300",
    x"01010100",
    x"10010001",
    x"0800A801",
    x"06010100",
    x"06020400",
    x"01020200",
    x"11000102",
    x"06020400",
    x"01020200",
    x"10020002",
    x"06010300",
    x"01010100",
    x"10010001",
    x"03010102",
    x"06020400",
    x"01020200",
    x"11000102",
    x"06010400",
    x"01010100",
    x"10010001",
    x"06020300",
    x"01020200",
    x"11000102",
    x"07008F00",
    x"07006900",
    x"07004300",
    x"06010000",
    x"01010100",
    x"10010001",
    x"0C000101",
    x"06010000",
    x"01010100",
    x"10010001",
    x"0C000101",
    x"06010200",
    x"06020200",
    x"01020200",
    x"11000102",
    x"06020200",
    x"01020200",
    x"10020002",
    x"06010000",
    x"01010100",
    x"10010001",
    x"02010102",
    x"06020200",
    x"01020200",
    x"11000102",
    x"06010200",
    x"01010100",
    x"10010001",
    x"06020000",
    x"01020200",
    x"11000102",
    x"07001100",
    OTHERS => (OTHERS => '0'));

    CONSTANT mem : mem_t := switch_chanel;
BEGIN
    data <= mem(conv_integer(addr));
END ARCHITECTURE;